module fmul (a, b, rm, s);
	input [31:0] a;		// fp a
	input [31:0] b;		// fp b
	input [1:0] rm;		// round mode
	output [31:0] s;	// fp output
	
	wire a_epxo_is_00 = ~|a[30:23];		// expo=00
	wire b_expo_is_00 = ~|b[30:23];
	wire a_expo_is_ff = &a[30:23];		// expo=ff
	wire b_expo_is_ff = &b[30:23];
	wire a_frac_is_00 = ~|a[22:0];		// frac=0
	wire b_frac_is_00 = ~|b[22:0];

	wire a_is_inf = a_expo_is_ff & a_frac_is_00;
	wire b_is_inf = b_expo_is_ff & b_frac_is_00;
	wire a_is_nan = a_expo_is_ff & ~a_frac_is_00;
	wire b_is_nan = b_expo_is_ff & ~b_frac_is_00;
	wire a_is_0 = a_expo_is_00 & a_frac_is_00;
	wire b_is_0 = b_expo_is_00 & b_frac_is_00;
	wire s_is_inf = a_is_inf | b_is_inf;
	wire s_is_nan = a_is_nan | b_is_nan | (a_is_inf&b_is_0) | (b_is_inf&a_is_0);
	
	wire [22:0] nan_frac = (a[21:0]>b[21:0])?{1'b1,a[21:0]}:{1'b1,b[21:0]};
	wire [22:0] inf_nan_frac = s_is_nan? nan_frac : 23'h0;
	
	wire sign = a[31]^b[31];
	wire [9:0] exp10 = {2'h0,a[30:23]} + {2'h0,b[30:23]} - 10'h7f + 
		a_expo_is_00 + b_expo_is_00;	// is a_expo is 00, expo10 add 1, so as b_expo is 0
	wire [23:0] a_frac24 = {~a_expo_is_00, a[22:0]};
	wire [23:0] b_frac24 = {~b_expo_is_00, b[22:0]};
	wire [47:0] z;
	wire [47:8] z_sum;
	wire [47:8] z_carry;

	// multiplication 1: carry and sum generated by wallace tree
	wallace_24x24 wt24 (a_frac24, b_frac24, z_sum, z_carry, z[7:0]);
	// multiplication 2: product by adding carry and sum
	assign z[47:8] = {1'b0, z_sum} + z_carry;	//xx.xxxxxxxx...
	// normalization
	wire [46:0] z5,z4,z3,z2,z1,z0;
	wire zero5,zero4,zero3,zero2,zero1,zero0;
	assign zero5 = ~|z[46:15];
	


endmodule
