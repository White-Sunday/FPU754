module pipelined_fadder (a,b,sub,rm,s,clk,clrn,e);
endmodule
